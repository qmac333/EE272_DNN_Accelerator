* Ring oscillator circuit

.subckt ringosc out vdd gnd

* YOUR IMPLEMENTATION HERE

.ends
