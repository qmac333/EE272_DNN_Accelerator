/home/users/jiajunc4/ee272/git_ee272/EE272_DNN_Accelerator/hw7/dnn-accelerator-pnr/ConvVerilog/build/3-skywater-130nm/view-standard/stdcells.lef