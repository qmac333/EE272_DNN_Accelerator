../../5-testbench/outputs/testbench.sv