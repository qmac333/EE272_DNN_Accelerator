* Testbench for a ring oscillator

* YOUR IMPLEMENTATION HERE

Vringosc V0 0 1.5
Vinv V1 0 1.8


Xringosc ro_out V0 0 ringosc
Xinverter ro_out out V1 0 inv1

* initialize ro_out to 0 to prevent the oscillator
* from starting the equilibrium point
.ic V(ro_out)=0

* specify simulation duration, with "uic"
* indicating "use initial conditions"
.tran 10e-12 25e-09 0e-00 uic

* ngspice control commands
* .control
* save all
* run
* write
* .endc

.control
let pwr=0.1
while pwr < 1.81
  set pwr = $&pwr
  alter V0 dc pwr
  save out
  run
  write sim_{$pwr}.raw out
  let pwr = pwr + 0.1
end
.endc

* end of the testbench
.end
