magic
tech sky130A
magscale 1 2
timestamp 1741243312
<< nwell >>
rect -101 271 2804 592
<< pwell >>
rect 29 -7 63 27
rect 444 -7 478 27
rect 859 -7 893 27
rect 1274 -7 1308 27
rect 1689 -7 1723 27
rect 2104 -7 2138 27
rect 2519 -7 2553 27
<< scnmos >>
rect 120 57 150 187
rect 535 57 565 187
rect 950 57 980 187
rect 1365 57 1395 187
rect 1780 57 1810 187
rect 2195 57 2225 187
rect 2610 57 2640 187
<< scpmoshvt >>
rect 120 307 150 507
rect 535 307 565 507
rect 950 307 980 507
rect 1365 307 1395 507
rect 1780 307 1810 507
rect 2195 307 2225 507
rect 2610 307 2640 507
<< ndiff >>
rect 68 175 120 187
rect 68 141 76 175
rect 110 141 120 175
rect 68 107 120 141
rect 68 73 76 107
rect 110 73 120 107
rect 68 57 120 73
rect 150 175 202 187
rect 150 141 160 175
rect 194 141 202 175
rect 150 107 202 141
rect 150 73 160 107
rect 194 73 202 107
rect 150 57 202 73
rect 483 175 535 187
rect 483 141 491 175
rect 525 141 535 175
rect 483 107 535 141
rect 483 73 491 107
rect 525 73 535 107
rect 483 57 535 73
rect 565 175 617 187
rect 565 141 575 175
rect 609 141 617 175
rect 565 107 617 141
rect 565 73 575 107
rect 609 73 617 107
rect 565 57 617 73
rect 898 175 950 187
rect 898 141 906 175
rect 940 141 950 175
rect 898 107 950 141
rect 898 73 906 107
rect 940 73 950 107
rect 898 57 950 73
rect 980 175 1032 187
rect 980 141 990 175
rect 1024 141 1032 175
rect 980 107 1032 141
rect 980 73 990 107
rect 1024 73 1032 107
rect 980 57 1032 73
rect 1313 175 1365 187
rect 1313 141 1321 175
rect 1355 141 1365 175
rect 1313 107 1365 141
rect 1313 73 1321 107
rect 1355 73 1365 107
rect 1313 57 1365 73
rect 1395 175 1447 187
rect 1395 141 1405 175
rect 1439 141 1447 175
rect 1395 107 1447 141
rect 1395 73 1405 107
rect 1439 73 1447 107
rect 1395 57 1447 73
rect 1728 175 1780 187
rect 1728 141 1736 175
rect 1770 141 1780 175
rect 1728 107 1780 141
rect 1728 73 1736 107
rect 1770 73 1780 107
rect 1728 57 1780 73
rect 1810 175 1862 187
rect 1810 141 1820 175
rect 1854 141 1862 175
rect 1810 107 1862 141
rect 1810 73 1820 107
rect 1854 73 1862 107
rect 1810 57 1862 73
rect 2143 175 2195 187
rect 2143 141 2151 175
rect 2185 141 2195 175
rect 2143 107 2195 141
rect 2143 73 2151 107
rect 2185 73 2195 107
rect 2143 57 2195 73
rect 2225 175 2277 187
rect 2225 141 2235 175
rect 2269 141 2277 175
rect 2225 107 2277 141
rect 2225 73 2235 107
rect 2269 73 2277 107
rect 2225 57 2277 73
rect 2558 175 2610 187
rect 2558 141 2566 175
rect 2600 141 2610 175
rect 2558 107 2610 141
rect 2558 73 2566 107
rect 2600 73 2610 107
rect 2558 57 2610 73
rect 2640 175 2692 187
rect 2640 141 2650 175
rect 2684 141 2692 175
rect 2640 107 2692 141
rect 2640 73 2650 107
rect 2684 73 2692 107
rect 2640 57 2692 73
<< pdiff >>
rect 68 495 120 507
rect 68 461 76 495
rect 110 461 120 495
rect 68 427 120 461
rect 68 393 76 427
rect 110 393 120 427
rect 68 359 120 393
rect 68 325 76 359
rect 110 325 120 359
rect 68 307 120 325
rect 150 495 202 507
rect 150 461 160 495
rect 194 461 202 495
rect 483 495 535 507
rect 150 427 202 461
rect 150 393 160 427
rect 194 393 202 427
rect 150 359 202 393
rect 150 325 160 359
rect 194 325 202 359
rect 483 461 491 495
rect 525 461 535 495
rect 483 427 535 461
rect 483 393 491 427
rect 525 393 535 427
rect 483 359 535 393
rect 150 307 202 325
rect 483 325 491 359
rect 525 325 535 359
rect 483 307 535 325
rect 565 495 617 507
rect 565 461 575 495
rect 609 461 617 495
rect 898 495 950 507
rect 565 427 617 461
rect 565 393 575 427
rect 609 393 617 427
rect 565 359 617 393
rect 565 325 575 359
rect 609 325 617 359
rect 898 461 906 495
rect 940 461 950 495
rect 898 427 950 461
rect 898 393 906 427
rect 940 393 950 427
rect 898 359 950 393
rect 565 307 617 325
rect 898 325 906 359
rect 940 325 950 359
rect 898 307 950 325
rect 980 495 1032 507
rect 980 461 990 495
rect 1024 461 1032 495
rect 1313 495 1365 507
rect 980 427 1032 461
rect 980 393 990 427
rect 1024 393 1032 427
rect 980 359 1032 393
rect 980 325 990 359
rect 1024 325 1032 359
rect 1313 461 1321 495
rect 1355 461 1365 495
rect 1313 427 1365 461
rect 1313 393 1321 427
rect 1355 393 1365 427
rect 1313 359 1365 393
rect 980 307 1032 325
rect 1313 325 1321 359
rect 1355 325 1365 359
rect 1313 307 1365 325
rect 1395 495 1447 507
rect 1395 461 1405 495
rect 1439 461 1447 495
rect 1728 495 1780 507
rect 1395 427 1447 461
rect 1395 393 1405 427
rect 1439 393 1447 427
rect 1395 359 1447 393
rect 1395 325 1405 359
rect 1439 325 1447 359
rect 1728 461 1736 495
rect 1770 461 1780 495
rect 1728 427 1780 461
rect 1728 393 1736 427
rect 1770 393 1780 427
rect 1728 359 1780 393
rect 1395 307 1447 325
rect 1728 325 1736 359
rect 1770 325 1780 359
rect 1728 307 1780 325
rect 1810 495 1862 507
rect 1810 461 1820 495
rect 1854 461 1862 495
rect 2143 495 2195 507
rect 1810 427 1862 461
rect 1810 393 1820 427
rect 1854 393 1862 427
rect 1810 359 1862 393
rect 1810 325 1820 359
rect 1854 325 1862 359
rect 2143 461 2151 495
rect 2185 461 2195 495
rect 2143 427 2195 461
rect 2143 393 2151 427
rect 2185 393 2195 427
rect 2143 359 2195 393
rect 1810 307 1862 325
rect 2143 325 2151 359
rect 2185 325 2195 359
rect 2143 307 2195 325
rect 2225 495 2277 507
rect 2225 461 2235 495
rect 2269 461 2277 495
rect 2558 495 2610 507
rect 2225 427 2277 461
rect 2225 393 2235 427
rect 2269 393 2277 427
rect 2225 359 2277 393
rect 2225 325 2235 359
rect 2269 325 2277 359
rect 2558 461 2566 495
rect 2600 461 2610 495
rect 2558 427 2610 461
rect 2558 393 2566 427
rect 2600 393 2610 427
rect 2558 359 2610 393
rect 2225 307 2277 325
rect 2558 325 2566 359
rect 2600 325 2610 359
rect 2558 307 2610 325
rect 2640 495 2692 507
rect 2640 461 2650 495
rect 2684 461 2692 495
rect 2640 427 2692 461
rect 2640 393 2650 427
rect 2684 393 2692 427
rect 2640 359 2692 393
rect 2640 325 2650 359
rect 2684 325 2692 359
rect 2640 307 2692 325
<< ndiffc >>
rect 76 141 110 175
rect 76 73 110 107
rect 160 141 194 175
rect 160 73 194 107
rect 491 141 525 175
rect 491 73 525 107
rect 575 141 609 175
rect 575 73 609 107
rect 906 141 940 175
rect 906 73 940 107
rect 990 141 1024 175
rect 990 73 1024 107
rect 1321 141 1355 175
rect 1321 73 1355 107
rect 1405 141 1439 175
rect 1405 73 1439 107
rect 1736 141 1770 175
rect 1736 73 1770 107
rect 1820 141 1854 175
rect 1820 73 1854 107
rect 2151 141 2185 175
rect 2151 73 2185 107
rect 2235 141 2269 175
rect 2235 73 2269 107
rect 2566 141 2600 175
rect 2566 73 2600 107
rect 2650 141 2684 175
rect 2650 73 2684 107
<< pdiffc >>
rect 76 461 110 495
rect 76 393 110 427
rect 76 325 110 359
rect 160 461 194 495
rect 160 393 194 427
rect 160 325 194 359
rect 491 461 525 495
rect 491 393 525 427
rect 491 325 525 359
rect 575 461 609 495
rect 575 393 609 427
rect 575 325 609 359
rect 906 461 940 495
rect 906 393 940 427
rect 906 325 940 359
rect 990 461 1024 495
rect 990 393 1024 427
rect 990 325 1024 359
rect 1321 461 1355 495
rect 1321 393 1355 427
rect 1321 325 1355 359
rect 1405 461 1439 495
rect 1405 393 1439 427
rect 1405 325 1439 359
rect 1736 461 1770 495
rect 1736 393 1770 427
rect 1736 325 1770 359
rect 1820 461 1854 495
rect 1820 393 1854 427
rect 1820 325 1854 359
rect 2151 461 2185 495
rect 2151 393 2185 427
rect 2151 325 2185 359
rect 2235 461 2269 495
rect 2235 393 2269 427
rect 2235 325 2269 359
rect 2566 461 2600 495
rect 2566 393 2600 427
rect 2566 325 2600 359
rect 2650 461 2684 495
rect 2650 393 2684 427
rect 2650 325 2684 359
<< psubdiff >>
rect -64 170 14 200
rect -64 91 -51 170
rect 1 91 14 170
rect -64 65 14 91
rect 351 170 429 200
rect 351 91 364 170
rect 416 91 429 170
rect 351 65 429 91
rect 766 170 844 200
rect 766 91 779 170
rect 831 91 844 170
rect 766 65 844 91
rect 1181 170 1259 200
rect 1181 91 1194 170
rect 1246 91 1259 170
rect 1181 65 1259 91
rect 1596 170 1674 200
rect 1596 91 1609 170
rect 1661 91 1674 170
rect 1596 65 1674 91
rect 2011 170 2089 200
rect 2011 91 2024 170
rect 2076 91 2089 170
rect 2011 65 2089 91
rect 2426 170 2504 200
rect 2426 91 2439 170
rect 2491 91 2504 170
rect 2426 65 2504 91
<< nsubdiff >>
rect -64 458 14 489
rect -64 395 -51 458
rect 3 395 14 458
rect -64 346 14 395
rect 351 458 429 489
rect 351 395 364 458
rect 418 395 429 458
rect 351 346 429 395
rect 766 458 844 489
rect 766 395 779 458
rect 833 395 844 458
rect 766 346 844 395
rect 1181 458 1259 489
rect 1181 395 1194 458
rect 1248 395 1259 458
rect 1181 346 1259 395
rect 1596 458 1674 489
rect 1596 395 1609 458
rect 1663 395 1674 458
rect 1596 346 1674 395
rect 2011 458 2089 489
rect 2011 395 2024 458
rect 2078 395 2089 458
rect 2011 346 2089 395
rect 2426 458 2504 489
rect 2426 395 2439 458
rect 2493 395 2504 458
rect 2426 346 2504 395
<< psubdiffcont >>
rect -51 91 1 170
rect 364 91 416 170
rect 779 91 831 170
rect 1194 91 1246 170
rect 1609 91 1661 170
rect 2024 91 2076 170
rect 2439 91 2491 170
<< nsubdiffcont >>
rect -51 395 3 458
rect 364 395 418 458
rect 779 395 833 458
rect 1194 395 1248 458
rect 1609 395 1663 458
rect 2024 395 2078 458
rect 2439 395 2493 458
<< poly >>
rect 120 507 150 533
rect 535 507 565 533
rect 950 507 980 533
rect 1365 507 1395 533
rect 1780 507 1810 533
rect 2195 507 2225 533
rect 2610 507 2640 533
rect 120 275 150 307
rect 535 275 565 307
rect 950 275 980 307
rect 1365 275 1395 307
rect 1780 275 1810 307
rect 2195 275 2225 307
rect 2610 275 2640 307
rect 64 259 150 275
rect 64 225 80 259
rect 114 225 150 259
rect 64 209 150 225
rect 479 259 565 275
rect 479 225 495 259
rect 529 225 565 259
rect 479 209 565 225
rect 894 259 980 275
rect 894 225 910 259
rect 944 225 980 259
rect 894 209 980 225
rect 1309 259 1395 275
rect 1309 225 1325 259
rect 1359 225 1395 259
rect 1309 209 1395 225
rect 1724 259 1810 275
rect 1724 225 1740 259
rect 1774 225 1810 259
rect 1724 209 1810 225
rect 2139 259 2225 275
rect 2139 225 2155 259
rect 2189 225 2225 259
rect 2139 209 2225 225
rect 2554 259 2640 275
rect 2554 225 2570 259
rect 2604 225 2640 259
rect 2554 209 2640 225
rect 120 187 150 209
rect 535 187 565 209
rect 950 187 980 209
rect 1365 187 1395 209
rect 1780 187 1810 209
rect 2195 187 2225 209
rect 2610 187 2640 209
rect 120 31 150 57
rect 535 31 565 57
rect 950 31 980 57
rect 1365 31 1395 57
rect 1780 31 1810 57
rect 2195 31 2225 57
rect 2610 31 2640 57
<< polycont >>
rect 80 225 114 259
rect 495 225 529 259
rect 910 225 944 259
rect 1325 225 1359 259
rect 1740 225 1774 259
rect 2155 225 2189 259
rect 2570 225 2604 259
<< locali >>
rect 0 537 29 571
rect 63 537 121 571
rect 155 537 213 571
rect 247 537 276 571
rect 415 537 444 571
rect 478 537 536 571
rect 570 537 628 571
rect 662 537 691 571
rect 830 537 859 571
rect 893 537 951 571
rect 985 537 1043 571
rect 1077 537 1106 571
rect 1245 537 1274 571
rect 1308 537 1366 571
rect 1400 537 1458 571
rect 1492 537 1521 571
rect 1660 537 1689 571
rect 1723 537 1781 571
rect 1815 537 1873 571
rect 1907 537 1936 571
rect 2075 537 2104 571
rect 2138 537 2196 571
rect 2230 537 2288 571
rect 2322 537 2351 571
rect 2490 537 2519 571
rect 2553 537 2611 571
rect 2645 537 2703 571
rect 2737 537 2766 571
rect 68 495 110 537
rect 68 476 76 495
rect -64 461 76 476
rect -64 458 110 461
rect -64 395 -51 458
rect 3 427 110 458
rect 3 395 76 427
rect -64 393 76 395
rect -64 369 110 393
rect 68 359 110 369
rect 68 325 76 359
rect 68 309 110 325
rect 144 495 210 503
rect 144 461 160 495
rect 194 461 210 495
rect 483 495 525 537
rect 483 476 491 495
rect 144 427 210 461
rect 144 393 160 427
rect 194 393 210 427
rect 144 359 210 393
rect 351 461 491 476
rect 351 458 525 461
rect 351 395 364 458
rect 418 427 525 458
rect 418 395 491 427
rect 351 393 491 395
rect 351 369 525 393
rect 144 325 160 359
rect 194 325 210 359
rect 144 307 210 325
rect 483 359 525 369
rect 483 325 491 359
rect 483 309 525 325
rect 559 495 625 503
rect 559 461 575 495
rect 609 461 625 495
rect 898 495 940 537
rect 898 476 906 495
rect 559 427 625 461
rect 559 393 575 427
rect 609 393 625 427
rect 559 359 625 393
rect 766 461 906 476
rect 766 458 940 461
rect 766 395 779 458
rect 833 427 940 458
rect 833 395 906 427
rect 766 393 906 395
rect 766 369 940 393
rect 559 325 575 359
rect 609 325 625 359
rect 559 307 625 325
rect 898 359 940 369
rect 898 325 906 359
rect 898 309 940 325
rect 974 495 1040 503
rect 974 461 990 495
rect 1024 461 1040 495
rect 1313 495 1355 537
rect 1313 476 1321 495
rect 974 427 1040 461
rect 974 393 990 427
rect 1024 393 1040 427
rect 974 359 1040 393
rect 1181 461 1321 476
rect 1181 458 1355 461
rect 1181 395 1194 458
rect 1248 427 1355 458
rect 1248 395 1321 427
rect 1181 393 1321 395
rect 1181 369 1355 393
rect 974 325 990 359
rect 1024 325 1040 359
rect 974 307 1040 325
rect 1313 359 1355 369
rect 1313 325 1321 359
rect 1313 309 1355 325
rect 1389 495 1455 503
rect 1389 461 1405 495
rect 1439 461 1455 495
rect 1728 495 1770 537
rect 1728 476 1736 495
rect 1389 427 1455 461
rect 1389 393 1405 427
rect 1439 393 1455 427
rect 1389 359 1455 393
rect 1596 461 1736 476
rect 1596 458 1770 461
rect 1596 395 1609 458
rect 1663 427 1770 458
rect 1663 395 1736 427
rect 1596 393 1736 395
rect 1596 369 1770 393
rect 1389 325 1405 359
rect 1439 325 1455 359
rect 1389 307 1455 325
rect 1728 359 1770 369
rect 1728 325 1736 359
rect 1728 309 1770 325
rect 1804 495 1870 503
rect 1804 461 1820 495
rect 1854 461 1870 495
rect 2143 495 2185 537
rect 2143 476 2151 495
rect 1804 427 1870 461
rect 1804 393 1820 427
rect 1854 393 1870 427
rect 1804 359 1870 393
rect 2011 461 2151 476
rect 2011 458 2185 461
rect 2011 395 2024 458
rect 2078 427 2185 458
rect 2078 395 2151 427
rect 2011 393 2151 395
rect 2011 369 2185 393
rect 1804 325 1820 359
rect 1854 325 1870 359
rect 1804 307 1870 325
rect 2143 359 2185 369
rect 2143 325 2151 359
rect 2143 309 2185 325
rect 2219 495 2285 503
rect 2219 461 2235 495
rect 2269 461 2285 495
rect 2558 495 2600 537
rect 2558 476 2566 495
rect 2219 427 2285 461
rect 2219 393 2235 427
rect 2269 393 2285 427
rect 2219 359 2285 393
rect 2426 461 2566 476
rect 2426 458 2600 461
rect 2426 395 2439 458
rect 2493 427 2600 458
rect 2493 395 2566 427
rect 2426 393 2566 395
rect 2426 369 2600 393
rect 2219 325 2235 359
rect 2269 325 2285 359
rect 2219 307 2285 325
rect 2558 359 2600 369
rect 2558 325 2566 359
rect 2558 309 2600 325
rect 2634 495 2700 503
rect 2634 461 2650 495
rect 2684 461 2700 495
rect 2634 427 2700 461
rect 2634 393 2650 427
rect 2684 393 2700 427
rect 2634 359 2700 393
rect 2634 325 2650 359
rect 2684 325 2700 359
rect 2634 307 2700 325
rect 164 273 210 307
rect 579 273 625 307
rect 994 273 1040 307
rect 1409 273 1455 307
rect 1824 273 1870 307
rect 2239 273 2285 307
rect 2654 273 2700 307
rect -239 259 130 273
rect -239 225 80 259
rect 114 225 130 259
rect 164 259 545 273
rect 164 225 495 259
rect 529 225 545 259
rect 579 259 960 273
rect 579 225 910 259
rect 944 225 960 259
rect 994 259 1375 273
rect 994 225 1325 259
rect 1359 225 1375 259
rect 1409 259 1790 273
rect 1409 225 1740 259
rect 1774 225 1790 259
rect 1824 259 2205 273
rect 1824 225 2155 259
rect 2189 225 2205 259
rect 2239 259 2620 273
rect 2239 225 2570 259
rect 2604 225 2620 259
rect 2654 225 2944 273
rect -239 -76 -191 225
rect -64 175 110 191
rect 164 187 210 225
rect -64 170 76 175
rect -64 91 -51 170
rect 1 141 76 170
rect 1 107 110 141
rect 1 91 76 107
rect -64 73 76 91
rect -64 72 110 73
rect 64 27 110 72
rect 144 175 210 187
rect 144 141 160 175
rect 194 141 210 175
rect 144 107 210 141
rect 144 73 160 107
rect 194 73 210 107
rect 144 61 210 73
rect 351 175 525 191
rect 579 187 625 225
rect 351 170 491 175
rect 351 91 364 170
rect 416 141 491 170
rect 416 107 525 141
rect 416 91 491 107
rect 351 73 491 91
rect 351 72 525 73
rect 479 27 525 72
rect 559 175 625 187
rect 559 141 575 175
rect 609 141 625 175
rect 559 107 625 141
rect 559 73 575 107
rect 609 73 625 107
rect 559 61 625 73
rect 766 175 940 191
rect 994 187 1040 225
rect 766 170 906 175
rect 766 91 779 170
rect 831 141 906 170
rect 831 107 940 141
rect 831 91 906 107
rect 766 73 906 91
rect 766 72 940 73
rect 894 27 940 72
rect 974 175 1040 187
rect 974 141 990 175
rect 1024 141 1040 175
rect 974 107 1040 141
rect 974 73 990 107
rect 1024 73 1040 107
rect 974 61 1040 73
rect 1181 175 1355 191
rect 1409 187 1455 225
rect 1181 170 1321 175
rect 1181 91 1194 170
rect 1246 141 1321 170
rect 1246 107 1355 141
rect 1246 91 1321 107
rect 1181 73 1321 91
rect 1181 72 1355 73
rect 1309 27 1355 72
rect 1389 175 1455 187
rect 1389 141 1405 175
rect 1439 141 1455 175
rect 1389 107 1455 141
rect 1389 73 1405 107
rect 1439 73 1455 107
rect 1389 61 1455 73
rect 1596 175 1770 191
rect 1824 187 1870 225
rect 1596 170 1736 175
rect 1596 91 1609 170
rect 1661 141 1736 170
rect 1661 107 1770 141
rect 1661 91 1736 107
rect 1596 73 1736 91
rect 1596 72 1770 73
rect 1724 27 1770 72
rect 1804 175 1870 187
rect 1804 141 1820 175
rect 1854 141 1870 175
rect 1804 107 1870 141
rect 1804 73 1820 107
rect 1854 73 1870 107
rect 1804 61 1870 73
rect 2011 175 2185 191
rect 2239 187 2285 225
rect 2011 170 2151 175
rect 2011 91 2024 170
rect 2076 141 2151 170
rect 2076 107 2185 141
rect 2076 91 2151 107
rect 2011 73 2151 91
rect 2011 72 2185 73
rect 2139 27 2185 72
rect 2219 175 2285 187
rect 2219 141 2235 175
rect 2269 141 2285 175
rect 2219 107 2285 141
rect 2219 73 2235 107
rect 2269 73 2285 107
rect 2219 61 2285 73
rect 2426 175 2600 191
rect 2654 187 2700 225
rect 2426 170 2566 175
rect 2426 91 2439 170
rect 2491 141 2566 170
rect 2491 107 2600 141
rect 2491 91 2566 107
rect 2426 73 2566 91
rect 2426 72 2600 73
rect 2554 27 2600 72
rect 2634 175 2700 187
rect 2634 141 2650 175
rect 2684 141 2700 175
rect 2634 107 2700 141
rect 2634 73 2650 107
rect 2684 73 2700 107
rect 2634 61 2700 73
rect 0 -7 29 27
rect 63 -7 121 27
rect 155 -7 213 27
rect 247 -7 276 27
rect 415 -7 444 27
rect 478 -7 536 27
rect 570 -7 628 27
rect 662 -7 691 27
rect 830 -7 859 27
rect 893 -7 951 27
rect 985 -7 1043 27
rect 1077 -7 1106 27
rect 1245 -7 1274 27
rect 1308 -7 1366 27
rect 1400 -7 1458 27
rect 1492 -7 1521 27
rect 1660 -7 1689 27
rect 1723 -7 1781 27
rect 1815 -7 1873 27
rect 1907 -7 1936 27
rect 2075 -7 2104 27
rect 2138 -7 2196 27
rect 2230 -7 2288 27
rect 2322 -7 2351 27
rect 2490 -7 2519 27
rect 2553 -7 2611 27
rect 2645 -7 2703 27
rect 2737 -7 2766 27
rect 2896 -76 2944 225
rect -239 -124 2944 -76
<< viali >>
rect 29 537 63 571
rect 121 537 155 571
rect 213 537 247 571
rect 444 537 478 571
rect 536 537 570 571
rect 628 537 662 571
rect 859 537 893 571
rect 951 537 985 571
rect 1043 537 1077 571
rect 1274 537 1308 571
rect 1366 537 1400 571
rect 1458 537 1492 571
rect 1689 537 1723 571
rect 1781 537 1815 571
rect 1873 537 1907 571
rect 2104 537 2138 571
rect 2196 537 2230 571
rect 2288 537 2322 571
rect 2519 537 2553 571
rect 2611 537 2645 571
rect 2703 537 2737 571
rect 29 -7 63 27
rect 121 -7 155 27
rect 213 -7 247 27
rect 444 -7 478 27
rect 536 -7 570 27
rect 628 -7 662 27
rect 859 -7 893 27
rect 951 -7 985 27
rect 1043 -7 1077 27
rect 1274 -7 1308 27
rect 1366 -7 1400 27
rect 1458 -7 1492 27
rect 1689 -7 1723 27
rect 1781 -7 1815 27
rect 1873 -7 1907 27
rect 2104 -7 2138 27
rect 2196 -7 2230 27
rect 2288 -7 2322 27
rect 2519 -7 2553 27
rect 2611 -7 2645 27
rect 2703 -7 2737 27
<< metal1 >>
rect -101 571 2804 602
rect -101 537 29 571
rect 63 537 121 571
rect 155 537 213 571
rect 247 537 444 571
rect 478 537 536 571
rect 570 537 628 571
rect 662 537 859 571
rect 893 537 951 571
rect 985 537 1043 571
rect 1077 537 1274 571
rect 1308 537 1366 571
rect 1400 537 1458 571
rect 1492 537 1689 571
rect 1723 537 1781 571
rect 1815 537 1873 571
rect 1907 537 2104 571
rect 2138 537 2196 571
rect 2230 537 2288 571
rect 2322 537 2519 571
rect 2553 537 2611 571
rect 2645 537 2703 571
rect 2737 537 2804 571
rect -101 506 2804 537
rect -101 27 2804 58
rect -101 -7 29 27
rect 63 -7 121 27
rect 155 -7 213 27
rect 247 -7 444 27
rect 478 -7 536 27
rect 570 -7 628 27
rect 662 -7 859 27
rect 893 -7 951 27
rect 985 -7 1043 27
rect 1077 -7 1274 27
rect 1308 -7 1366 27
rect 1400 -7 1458 27
rect 1492 -7 1689 27
rect 1723 -7 1781 27
rect 1815 -7 1873 27
rect 1907 -7 2104 27
rect 2138 -7 2196 27
rect 2230 -7 2288 27
rect 2322 -7 2519 27
rect 2553 -7 2611 27
rect 2645 -7 2703 27
rect 2737 -7 2804 27
rect -101 -38 2804 -7
<< labels >>
flabel locali 2716 230 2759 267 1 FreeSans 400 0 0 0 out
port 1 n
flabel metal1 1548 -9 1598 28 1 FreeSans 400 0 0 0 gnd
port 3 n
flabel locali 72 231 106 265 0 FreeSans 340 0 0 0 inv1_0[0].A
flabel locali 164 299 198 333 0 FreeSans 340 0 0 0 inv1_0[0].Y
flabel metal1 29 537 63 571 0 FreeSans 200 0 0 0 inv1_0[0].VPWR
flabel metal1 29 -7 63 27 0 FreeSans 200 0 0 0 inv1_0[0].VGND
rlabel comment 0 10 0 10 4 inv1_0[0].inv_1
flabel locali 487 231 521 265 0 FreeSans 340 0 0 0 inv1_0[1].A
flabel locali 579 299 613 333 0 FreeSans 340 0 0 0 inv1_0[1].Y
flabel metal1 444 537 478 571 0 FreeSans 200 0 0 0 inv1_0[1].VPWR
flabel metal1 444 -7 478 27 0 FreeSans 200 0 0 0 inv1_0[1].VGND
rlabel comment 415 10 415 10 4 inv1_0[1].inv_1
flabel locali 902 231 936 265 0 FreeSans 340 0 0 0 inv1_0[2].A
flabel locali 994 299 1028 333 0 FreeSans 340 0 0 0 inv1_0[2].Y
flabel metal1 859 537 893 571 0 FreeSans 200 0 0 0 inv1_0[2].VPWR
flabel metal1 859 -7 893 27 0 FreeSans 200 0 0 0 inv1_0[2].VGND
rlabel comment 830 10 830 10 4 inv1_0[2].inv_1
flabel locali 1317 231 1351 265 0 FreeSans 340 0 0 0 inv1_0[3].A
flabel locali 1409 299 1443 333 0 FreeSans 340 0 0 0 inv1_0[3].Y
flabel metal1 1274 537 1308 571 0 FreeSans 200 0 0 0 inv1_0[3].VPWR
flabel metal1 1274 -7 1308 27 0 FreeSans 200 0 0 0 inv1_0[3].VGND
rlabel comment 1245 10 1245 10 4 inv1_0[3].inv_1
flabel locali 1732 231 1766 265 0 FreeSans 340 0 0 0 inv1_0[4].A
flabel locali 1824 299 1858 333 0 FreeSans 340 0 0 0 inv1_0[4].Y
flabel metal1 1689 537 1723 571 0 FreeSans 200 0 0 0 inv1_0[4].VPWR
flabel metal1 1689 -7 1723 27 0 FreeSans 200 0 0 0 inv1_0[4].VGND
rlabel comment 1660 10 1660 10 4 inv1_0[4].inv_1
flabel locali 2147 231 2181 265 0 FreeSans 340 0 0 0 inv1_0[5].A
flabel locali 2239 299 2273 333 0 FreeSans 340 0 0 0 inv1_0[5].Y
flabel metal1 2104 537 2138 571 0 FreeSans 200 0 0 0 inv1_0[5].VPWR
flabel metal1 2104 -7 2138 27 0 FreeSans 200 0 0 0 inv1_0[5].VGND
rlabel comment 2075 10 2075 10 4 inv1_0[5].inv_1
flabel locali 2562 231 2596 265 0 FreeSans 340 0 0 0 inv1_0[6].A
flabel locali 2654 299 2688 333 0 FreeSans 340 0 0 0 inv1_0[6].Y
flabel metal1 2519 537 2553 571 0 FreeSans 200 0 0 0 inv1_0[6].VPWR
flabel metal1 2519 -7 2553 27 0 FreeSans 200 0 0 0 inv1_0[6].VGND
rlabel comment 2490 10 2490 10 4 inv1_0[6].inv_1
flabel metal1 1536 537 1588 576 1 FreeSans 400 0 0 0 vdd
port 2 n
<< end >>
