VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MACRO sky130_sram_1kbyte_1rw1r_32x256_8
   CLASS BLOCK ;
   SIZE 481.14 BY 400.22 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  107.44 0.0 107.82 1.06 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  113.56 0.0 113.94 1.06 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  119.0 0.0 119.38 1.06 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  125.8 0.0 126.18 1.06 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  131.24 0.0 131.62 1.06 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  136.68 0.0 137.06 1.06 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  142.12 0.0 142.5 1.06 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  148.92 0.0 149.3 1.06 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  154.36 0.0 154.74 1.06 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  159.8 0.0 160.18 1.06 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  165.92 0.0 166.3 1.06 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  171.36 0.0 171.74 1.06 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  178.16 0.0 178.54 1.06 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  183.6 0.0 183.98 1.06 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  189.04 0.0 189.42 1.06 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  195.16 0.0 195.54 1.06 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  201.96 0.0 202.34 1.06 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  207.4 0.0 207.78 1.06 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  212.84 0.0 213.22 1.06 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  218.28 0.0 218.66 1.06 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  225.08 0.0 225.46 1.06 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  230.52 0.0 230.9 1.06 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  235.96 0.0 236.34 1.06 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  242.08 0.0 242.46 1.06 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  247.52 0.0 247.9 1.06 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  254.32 0.0 254.7 1.06 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  259.76 0.0 260.14 1.06 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  265.2 0.0 265.58 1.06 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  270.64 0.0 271.02 1.06 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  276.76 0.0 277.14 1.06 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  283.56 0.0 283.94 1.06 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  289.0 0.0 289.38 1.06 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  78.2 0.0 78.58 1.06 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 129.88 1.06 130.26 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 138.04 1.06 138.42 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 143.48 1.06 143.86 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 151.64 1.06 152.02 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 157.08 1.06 157.46 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 165.92 1.06 166.3 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 171.36 1.06 171.74 ;
      END
   END addr0[7]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  397.8 399.16 398.18 400.22 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  480.08 84.32 481.14 84.7 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  480.08 76.16 481.14 76.54 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  480.08 70.72 481.14 71.1 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  416.16 0.0 416.54 1.06 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  414.12 0.0 414.5 1.06 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  414.8 0.0 415.18 1.06 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  415.48 0.0 415.86 1.06 ;
      END
   END addr1[7]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 28.56 1.06 28.94 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  480.08 383.52 481.14 383.9 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 36.72 1.06 37.1 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  29.92 0.0 30.3 1.06 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  450.84 399.16 451.22 400.22 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  84.32 0.0 84.7 1.06 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  89.76 0.0 90.14 1.06 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  96.56 0.0 96.94 1.06 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  101.32 0.0 101.7 1.06 ;
      END
   END wmask0[3]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  140.08 0.0 140.46 1.06 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  146.88 0.0 147.26 1.06 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  152.32 0.0 152.7 1.06 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  160.48 0.0 160.86 1.06 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  166.6 0.0 166.98 1.06 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.72 0.0 173.1 1.06 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.84 0.0 179.22 1.06 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  184.96 0.0 185.34 1.06 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  189.72 0.0 190.1 1.06 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.2 0.0 197.58 1.06 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  204.0 0.0 204.38 1.06 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  210.12 0.0 210.5 1.06 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  216.24 0.0 216.62 1.06 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  222.36 0.0 222.74 1.06 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  228.48 0.0 228.86 1.06 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  233.92 0.0 234.3 1.06 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  240.04 0.0 240.42 1.06 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  246.16 0.0 246.54 1.06 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  253.64 0.0 254.02 1.06 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  257.72 0.0 258.1 1.06 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  266.56 0.0 266.94 1.06 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  272.68 0.0 273.06 1.06 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  278.8 0.0 279.18 1.06 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  284.92 0.0 285.3 1.06 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  289.68 0.0 290.06 1.06 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  297.16 0.0 297.54 1.06 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  303.28 0.0 303.66 1.06 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  310.08 0.0 310.46 1.06 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  316.2 0.0 316.58 1.06 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  322.32 0.0 322.7 1.06 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  328.44 0.0 328.82 1.06 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  334.56 0.0 334.94 1.06 ;
      END
   END dout0[31]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  141.44 399.16 141.82 400.22 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  148.24 399.16 148.62 400.22 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  153.68 399.16 154.06 400.22 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  160.48 399.16 160.86 400.22 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  166.6 399.16 166.98 400.22 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  173.4 399.16 173.78 400.22 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  179.52 399.16 179.9 400.22 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  184.96 399.16 185.34 400.22 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  191.76 399.16 192.14 400.22 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.2 399.16 197.58 400.22 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  204.0 399.16 204.38 400.22 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  210.12 399.16 210.5 400.22 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  216.92 399.16 217.3 400.22 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  222.36 399.16 222.74 400.22 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  228.48 399.16 228.86 400.22 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  235.28 399.16 235.66 400.22 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  241.4 399.16 241.78 400.22 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  248.2 399.16 248.58 400.22 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  253.64 399.16 254.02 400.22 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  260.44 399.16 260.82 400.22 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  265.88 399.16 266.26 400.22 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  272.0 399.16 272.38 400.22 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  278.8 399.16 279.18 400.22 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  284.92 399.16 285.3 400.22 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  291.72 399.16 292.1 400.22 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  297.16 399.16 297.54 400.22 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  303.96 399.16 304.34 400.22 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  310.08 399.16 310.46 400.22 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  316.88 399.16 317.26 400.22 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  322.32 399.16 322.7 400.22 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  328.44 399.16 328.82 400.22 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  335.24 399.16 335.62 400.22 ;
      END
   END dout1[31]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  4.76 4.76 6.5 395.46 ;
         LAYER met4 ;
         RECT  474.64 4.76 476.38 395.46 ;
         LAYER met3 ;
         RECT  4.76 393.72 476.38 395.46 ;
         LAYER met3 ;
         RECT  4.76 4.76 476.38 6.5 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  478.04 1.36 479.78 398.86 ;
         LAYER met3 ;
         RECT  1.36 397.12 479.78 398.86 ;
         LAYER met4 ;
         RECT  1.36 1.36 3.1 398.86 ;
         LAYER met3 ;
         RECT  1.36 1.36 479.78 3.1 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 480.52 399.6 ;
   LAYER  met2 ;
      RECT  0.62 0.62 480.52 399.6 ;
   LAYER  met3 ;
      RECT  1.66 129.28 480.52 130.86 ;
      RECT  0.62 130.86 1.66 137.44 ;
      RECT  0.62 139.02 1.66 142.88 ;
      RECT  0.62 144.46 1.66 151.04 ;
      RECT  0.62 152.62 1.66 156.48 ;
      RECT  0.62 158.06 1.66 165.32 ;
      RECT  0.62 166.9 1.66 170.76 ;
      RECT  1.66 83.72 479.48 85.3 ;
      RECT  1.66 85.3 479.48 129.28 ;
      RECT  479.48 85.3 480.52 129.28 ;
      RECT  479.48 77.14 480.52 83.72 ;
      RECT  479.48 71.7 480.52 75.56 ;
      RECT  1.66 130.86 479.48 382.92 ;
      RECT  1.66 382.92 479.48 384.5 ;
      RECT  479.48 130.86 480.52 382.92 ;
      RECT  0.62 29.54 1.66 36.12 ;
      RECT  0.62 37.7 1.66 129.28 ;
      RECT  1.66 384.5 4.16 393.12 ;
      RECT  1.66 393.12 4.16 396.06 ;
      RECT  4.16 384.5 476.98 393.12 ;
      RECT  476.98 384.5 479.48 393.12 ;
      RECT  476.98 393.12 479.48 396.06 ;
      RECT  1.66 4.16 4.16 7.1 ;
      RECT  1.66 7.1 4.16 83.72 ;
      RECT  4.16 7.1 476.98 83.72 ;
      RECT  476.98 4.16 479.48 7.1 ;
      RECT  476.98 7.1 479.48 83.72 ;
      RECT  0.62 172.34 0.76 396.52 ;
      RECT  0.62 396.52 0.76 399.46 ;
      RECT  0.62 399.46 0.76 399.6 ;
      RECT  0.76 172.34 1.66 396.52 ;
      RECT  0.76 399.46 1.66 399.6 ;
      RECT  479.48 384.5 480.38 396.52 ;
      RECT  479.48 399.46 480.38 399.6 ;
      RECT  480.38 384.5 480.52 396.52 ;
      RECT  480.38 396.52 480.52 399.46 ;
      RECT  480.38 399.46 480.52 399.6 ;
      RECT  1.66 396.06 4.16 396.52 ;
      RECT  1.66 399.46 4.16 399.6 ;
      RECT  4.16 396.06 476.98 396.52 ;
      RECT  4.16 399.46 476.98 399.6 ;
      RECT  476.98 396.06 479.48 396.52 ;
      RECT  476.98 399.46 479.48 399.6 ;
      RECT  479.48 0.62 480.38 0.76 ;
      RECT  479.48 3.7 480.38 70.12 ;
      RECT  480.38 0.62 480.52 0.76 ;
      RECT  480.38 0.76 480.52 3.7 ;
      RECT  480.38 3.7 480.52 70.12 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 3.7 ;
      RECT  0.62 3.7 0.76 27.96 ;
      RECT  0.76 0.62 1.66 0.76 ;
      RECT  0.76 3.7 1.66 27.96 ;
      RECT  1.66 0.62 4.16 0.76 ;
      RECT  1.66 3.7 4.16 4.16 ;
      RECT  4.16 0.62 476.98 0.76 ;
      RECT  4.16 3.7 476.98 4.16 ;
      RECT  476.98 0.62 479.48 0.76 ;
      RECT  476.98 3.7 479.48 4.16 ;
   LAYER  met4 ;
      RECT  106.84 1.66 108.42 399.6 ;
      RECT  108.42 0.62 112.96 1.66 ;
      RECT  114.54 0.62 118.4 1.66 ;
      RECT  119.98 0.62 125.2 1.66 ;
      RECT  126.78 0.62 130.64 1.66 ;
      RECT  132.22 0.62 136.08 1.66 ;
      RECT  155.34 0.62 159.2 1.66 ;
      RECT  260.74 0.62 264.6 1.66 ;
      RECT  108.42 1.66 397.2 398.56 ;
      RECT  397.2 1.66 398.78 398.56 ;
      RECT  30.9 0.62 77.6 1.66 ;
      RECT  398.78 398.56 450.24 399.6 ;
      RECT  79.18 0.62 83.72 1.66 ;
      RECT  85.3 0.62 89.16 1.66 ;
      RECT  90.74 0.62 95.96 1.66 ;
      RECT  97.54 0.62 100.72 1.66 ;
      RECT  102.3 0.62 106.84 1.66 ;
      RECT  137.66 0.62 139.48 1.66 ;
      RECT  141.06 0.62 141.52 1.66 ;
      RECT  143.1 0.62 146.28 1.66 ;
      RECT  147.86 0.62 148.32 1.66 ;
      RECT  149.9 0.62 151.72 1.66 ;
      RECT  153.3 0.62 153.76 1.66 ;
      RECT  161.46 0.62 165.32 1.66 ;
      RECT  167.58 0.62 170.76 1.66 ;
      RECT  173.7 0.62 177.56 1.66 ;
      RECT  179.82 0.62 183.0 1.66 ;
      RECT  185.94 0.62 188.44 1.66 ;
      RECT  190.7 0.62 194.56 1.66 ;
      RECT  196.14 0.62 196.6 1.66 ;
      RECT  198.18 0.62 201.36 1.66 ;
      RECT  202.94 0.62 203.4 1.66 ;
      RECT  204.98 0.62 206.8 1.66 ;
      RECT  208.38 0.62 209.52 1.66 ;
      RECT  211.1 0.62 212.24 1.66 ;
      RECT  213.82 0.62 215.64 1.66 ;
      RECT  217.22 0.62 217.68 1.66 ;
      RECT  219.26 0.62 221.76 1.66 ;
      RECT  223.34 0.62 224.48 1.66 ;
      RECT  226.06 0.62 227.88 1.66 ;
      RECT  229.46 0.62 229.92 1.66 ;
      RECT  231.5 0.62 233.32 1.66 ;
      RECT  234.9 0.62 235.36 1.66 ;
      RECT  236.94 0.62 239.44 1.66 ;
      RECT  241.02 0.62 241.48 1.66 ;
      RECT  243.06 0.62 245.56 1.66 ;
      RECT  248.5 0.62 253.04 1.66 ;
      RECT  255.3 0.62 257.12 1.66 ;
      RECT  258.7 0.62 259.16 1.66 ;
      RECT  267.54 0.62 270.04 1.66 ;
      RECT  271.62 0.62 272.08 1.66 ;
      RECT  273.66 0.62 276.16 1.66 ;
      RECT  277.74 0.62 278.2 1.66 ;
      RECT  279.78 0.62 282.96 1.66 ;
      RECT  285.9 0.62 288.4 1.66 ;
      RECT  290.66 0.62 296.56 1.66 ;
      RECT  298.14 0.62 302.68 1.66 ;
      RECT  304.26 0.62 309.48 1.66 ;
      RECT  311.06 0.62 315.6 1.66 ;
      RECT  317.18 0.62 321.72 1.66 ;
      RECT  323.3 0.62 327.84 1.66 ;
      RECT  329.42 0.62 333.96 1.66 ;
      RECT  335.54 0.62 413.52 1.66 ;
      RECT  108.42 398.56 140.84 399.6 ;
      RECT  142.42 398.56 147.64 399.6 ;
      RECT  149.22 398.56 153.08 399.6 ;
      RECT  154.66 398.56 159.88 399.6 ;
      RECT  161.46 398.56 166.0 399.6 ;
      RECT  167.58 398.56 172.8 399.6 ;
      RECT  174.38 398.56 178.92 399.6 ;
      RECT  180.5 398.56 184.36 399.6 ;
      RECT  185.94 398.56 191.16 399.6 ;
      RECT  192.74 398.56 196.6 399.6 ;
      RECT  198.18 398.56 203.4 399.6 ;
      RECT  204.98 398.56 209.52 399.6 ;
      RECT  211.1 398.56 216.32 399.6 ;
      RECT  217.9 398.56 221.76 399.6 ;
      RECT  223.34 398.56 227.88 399.6 ;
      RECT  229.46 398.56 234.68 399.6 ;
      RECT  236.26 398.56 240.8 399.6 ;
      RECT  242.38 398.56 247.6 399.6 ;
      RECT  249.18 398.56 253.04 399.6 ;
      RECT  254.62 398.56 259.84 399.6 ;
      RECT  261.42 398.56 265.28 399.6 ;
      RECT  266.86 398.56 271.4 399.6 ;
      RECT  272.98 398.56 278.2 399.6 ;
      RECT  279.78 398.56 284.32 399.6 ;
      RECT  285.9 398.56 291.12 399.6 ;
      RECT  292.7 398.56 296.56 399.6 ;
      RECT  298.14 398.56 303.36 399.6 ;
      RECT  304.94 398.56 309.48 399.6 ;
      RECT  311.06 398.56 316.28 399.6 ;
      RECT  317.86 398.56 321.72 399.6 ;
      RECT  323.3 398.56 327.84 399.6 ;
      RECT  329.42 398.56 334.64 399.6 ;
      RECT  336.22 398.56 397.2 399.6 ;
      RECT  4.16 1.66 7.1 4.16 ;
      RECT  4.16 396.06 7.1 399.6 ;
      RECT  7.1 1.66 106.84 4.16 ;
      RECT  7.1 4.16 106.84 396.06 ;
      RECT  7.1 396.06 106.84 399.6 ;
      RECT  398.78 1.66 474.04 4.16 ;
      RECT  398.78 4.16 474.04 396.06 ;
      RECT  398.78 396.06 474.04 398.56 ;
      RECT  474.04 1.66 476.98 4.16 ;
      RECT  474.04 396.06 476.98 398.56 ;
      RECT  417.14 0.62 477.44 0.76 ;
      RECT  417.14 0.76 477.44 1.66 ;
      RECT  477.44 0.62 480.38 0.76 ;
      RECT  480.38 0.62 480.52 0.76 ;
      RECT  480.38 0.76 480.52 1.66 ;
      RECT  451.82 398.56 477.44 399.46 ;
      RECT  451.82 399.46 477.44 399.6 ;
      RECT  477.44 399.46 480.38 399.6 ;
      RECT  480.38 398.56 480.52 399.46 ;
      RECT  480.38 399.46 480.52 399.6 ;
      RECT  476.98 1.66 477.44 4.16 ;
      RECT  480.38 1.66 480.52 4.16 ;
      RECT  476.98 4.16 477.44 396.06 ;
      RECT  480.38 4.16 480.52 396.06 ;
      RECT  476.98 396.06 477.44 398.56 ;
      RECT  480.38 396.06 480.52 398.56 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 1.66 ;
      RECT  0.76 0.62 3.7 0.76 ;
      RECT  3.7 0.62 29.32 0.76 ;
      RECT  3.7 0.76 29.32 1.66 ;
      RECT  0.62 1.66 0.76 4.16 ;
      RECT  3.7 1.66 4.16 4.16 ;
      RECT  0.62 4.16 0.76 396.06 ;
      RECT  3.7 4.16 4.16 396.06 ;
      RECT  0.62 396.06 0.76 399.46 ;
      RECT  0.62 399.46 0.76 399.6 ;
      RECT  0.76 399.46 3.7 399.6 ;
      RECT  3.7 396.06 4.16 399.46 ;
      RECT  3.7 399.46 4.16 399.6 ;
   END
END    sky130_sram_1kbyte_1rw1r_32x256_8
END    LIBRARY
