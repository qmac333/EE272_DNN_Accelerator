* Testbench for a ring oscillator

* YOUR IMPLEMENTATION HERE

* .param V0_sthelse 

Vringosc V0 0 1.5
Vinv V1 0 1.8


Xringosc ro_out V0 0 ringosc
Xinverter ro_out out V1 0 inv1

* initialize ro_out to 0 to prevent the oscillator
* from starting the equilibrium point
.ic V(ro_out)=0

* specify simulation duration, with "uic"
* indicating "use initial conditions"
.tran 10e-12 25e-09 0e-00 uic

* ngspice control commands
* .control
* save all
* run
* write
* .endc

.control
let pwr=0.1
while pwr < 1.81
  set pwr = $&pwr
  alter Vringosc dc pwr
  save out
  run
  write sim_{$pwr}.raw out
  let pwr = pwr + 0.1
  meas tran t_osc TRIG v(out) val=0.9 rise=2 TARG v(out) val=0.9 rise=3
end
.endc

* .meas tran t_osc TRIG v(out) val=0.9 rise=2 TARG v(out) val=0.9 rise=3

* end of the testbench
.end
