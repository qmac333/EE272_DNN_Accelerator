/home/users/jiajunc4/ee272/git_ee272/EE272_DNN_Accelerator/hw7/dnn-accelerator-pnr/ConvVerilog/build/4-sram/outputs/sky130_sram_4kbyte_1rw1r_32x1024_8.lef